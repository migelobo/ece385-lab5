module reg_file(
	input logic  [15:0] bus_data,
	input logic  [2:0] DRMUX_result,SR1MUX_result, lower3_SR2,
	input logic  LD_REG,
	output logic [15:0] SR2_OUT, SR1_OUT
);

logic [15:0] register[7:0];


endmodule 